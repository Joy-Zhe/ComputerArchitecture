`timescale 1ns / 1ps

module Bin2BCD(
    input [4:0]Binary,
    output [7:0]BCD
);

    //  HEX0-31  ===>   BCD编码
    
    wire x00 = Binary == 5'b00000;  //  00
    wire x01 = Binary == 5'b00001;  //  01
    wire x02 = Binary == 5'b00010;  //  02
    wire x03 = Binary == 5'b00011;  //  03
    wire x04 = Binary == 5'b00100;  //  04
    wire x05 = Binary == 5'b00101;  //  05
    wire x06 = Binary == 5'b00110;  //  06
    wire x07 = Binary == 5'b00111;  //  07

    wire x08 = Binary == 5'b01000;  //  08
    wire x09 = Binary == 5'b01001;  //  09
    wire x10 = Binary == 5'b01010;  //  10
    wire x11 = Binary == 5'b01011;  //  11
    wire x12 = Binary == 5'b01100;  //  12
    wire x13 = Binary == 5'b01101;  //  13
    wire x14 = Binary == 5'b01110;  //  14
    wire x15 = Binary == 5'b01111;  //  15

    wire x16 = Binary == 5'b10000;  //  16
    wire x17 = Binary == 5'b10001;  //  17
    wire x18 = Binary == 5'b10010;  //  18
    wire x19 = Binary == 5'b10011;  //  19
    wire x20 = Binary == 5'b10100;  //  20
    wire x21 = Binary == 5'b10101;  //  21
    wire x22 = Binary == 5'b10110;  //  22
    wire x23 = Binary == 5'b10111;  //  23

    wire x24 = Binary == 5'b11000;  //  24
    wire x25 = Binary == 5'b11001;  //  25
    wire x26 = Binary == 5'b11010;  //  26
    wire x27 = Binary == 5'b11011;  //  27
    wire x28 = Binary == 5'b11100;  //  28
    wire x29 = Binary == 5'b11101;  //  29
    wire x30 = Binary == 5'b11110;  //  30
    wire x31 = Binary == 5'b11111;  //  31
        
    assign BCD =    { {8{x00}}  &   8'b0000_0000 }   |  //  00
                    { {8{x01}}  &   8'b0000_0001 }   |  //  01
                    { {8{x02}}  &   8'b0000_0010 }   |  //  02
                    { {8{x03}}  &   8'b0000_0011 }   |  //  03
                    { {8{x04}}  &   8'b0000_0100 }   |  //  04
                    { {8{x05}}  &   8'b0000_0101 }   |  //  05
                    { {8{x06}}  &   8'b0000_0110 }   |  //  06
                    { {8{x07}}  &   8'b0000_0111 }   |  //  07

                    { {8{x08}}  &   8'b0000_1000 }   |  //  08
                    { {8{x09}}  &   8'b0000_1001 }   |  //  09
                    { {8{x10}}  &   8'b0001_0000 }   |  //  10
                    { {8{x11}}  &   8'b0001_0001 }   |  //  11
                    { {8{x12}}  &   8'b0001_0010 }   |  //  12
                    { {8{x13}}  &   8'b0001_0011 }   |  //  13
                    { {8{x14}}  &   8'b0001_0100 }   |  //  14
                    { {8{x15}}  &   8'b0001_0101 }   |  //  15

                    { {8{x16}}  &   8'b0001_0110 }   |  //  16
                    { {8{x17}}  &   8'b0001_0111 }   |  //  17
                    { {8{x18}}  &   8'b0001_1000 }   |  //  18
                    { {8{x19}}  &   8'b0001_1001 }   |  //  19
                    { {8{x20}}  &   8'b0010_0000 }   |  //  20
                    { {8{x21}}  &   8'b0010_0001 }   |  //  21
                    { {8{x22}}  &   8'b0010_0010 }   |  //  22
                    { {8{x23}}  &   8'b0010_0011 }   |  //  23

                    { {8{x24}}  &   8'b0010_0100 }   |  //  24
                    { {8{x25}}  &   8'b0010_0101 }   |  //  25
                    { {8{x26}}  &   8'b0010_0110 }   |  //  26
                    { {8{x27}}  &   8'b0010_0111 }   |  //  27
                    { {8{x28}}  &   8'b0010_1000 }   |  //  28
                    { {8{x29}}  &   8'b0010_1001 }   |  //  29
                    { {8{x30}}  &   8'b0011_0000 }   |  //  30
                    { {8{x31}}  &   8'b0011_0001 }   ;  //  31

    
endmodule
